module or_4_bit (
    input wire a,
    input wire b,
    input wire c,
    input wire d,
    output wire s  
);

assign s = a || b || c || d;


endmodule