`include "SSBR_4_bits/SSBR_4_bits.v"

module FIFO_8_4 (
    input wire clk,
    input wire D
);

SSBR_4_bits SSBR_4_bits_0();

endmodule