`include "SSBR_4_bits/SSBR_4_bits.v"

module LIFO_8_4.v (
    input wire clock,
    input wire D,

);




    
endmodule