module and_1_bit (
    input wire a0,
    input wire a1,
    output wire s
);

assign s = a0 & a1;
    
endmodule